module light(
	input  clk,
	input  rst,
	input  ps2_clk,
	input  ps2_data,
	
	output [7:0] data,
	input  allowin,  
	output data_valid

);
endmodule
