module mem1(
  input   clock,
  input   reset
);
  d_mem Memory ( // @[src/src/memory/Mem.scala 20:28]
  );
endmodule
